// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "ibex_xif_icache_core_base_seq.sv"
`include "ibex_xif_icache_core_back_line_seq.sv"
